�� sr piggeon.engine.SaveState�V v��� L stagest Ljava/util/HashMap;xpsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      sr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   sr test.ExampleStage�6H�ѫi  xr piggeon.engine.Stage�4�)�JOJ L camerat Lpiggeon/engine/Camera;L rootNodet Lpiggeon/engine/Node;L 
updateListt Ljava/util/LinkedList;xpsr piggeon.engine.Camera�QL-L� L 
cameraNodeq ~ xpsr piggeon.engine.Node(L��K��\ F rotationF scaleXF scaleYF xF yL childrent Ljava/util/ArrayList;L nodeNamet Ljava/lang/String;xp    ?�  ?�          sr java.util.ArrayListx����a� I sizexp   w   sr test.ExampleMovingBoxObject.�yս� J aI delaybI delayxI dxI dyxr piggeon.engine.GameObjectWv���y F heightI 	textureIDI vaoIDF widthL animatort Lpiggeon/engine/Animator;L goUpdatablesq ~ xq ~     ?�  ?�  C� CA  sq ~     w    xt  BH        BH  sr piggeon.engine.Animator�镳q&�� I currentFrameIndexI currentSpriteIndexZ loopingL idq ~ L spriteTimeTableq ~ L targetGameObjectt Lpiggeon/engine/GameObject;xp       t 	box_colorsq ~    w   ur [Ljava.lang.Object;��X�s)l  xp   sr piggeon.util.ImageInfo���B�0 I heightI 	textureIDI widthxp   2      2sq ~    uq ~ !   sq ~ #   2      2q ~ %uq ~ !   sq ~ #   2      2q ~ %uq ~ !   sq ~ #   2      2q ~ %xq ~ sq ~     w    x      �           ����sr test.TextBoxExampleObject�L"��P J xL infot Lpiggeon/util/ImageInfo;xq ~     ?�  ?�  Cz  Cz  sq ~     w    xq ~ B�        B�  psq ~     w    x        sq ~ #   x      xxq ~ q ~ sr java.util.LinkedList)S]J`�"  xpw   q ~ q ~ /sr test.SoundExampleObject0��p�=�� J cdxq ~     ?�  ?�          sq ~     w    xq ~                 psq ~     w    x      1xx